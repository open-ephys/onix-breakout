// NB: colors.mem was generated using colors.py. There are lots of hardcoded
// constants in here that would need to be changed if the number of colors or
// their order is altered

`include "./ws2811/ws2811.v"

module neopix_controller # (
    parameter CLK_RATE_HZ = 50_000_000
) (
    // Clock and reset
    input   wire            i_clk,
    input   wire            i_reset,

    // Derived from host to breakout slow word
    input   wire            i_acq_running,
    input   wire            i_acq_reset_done,
    input   wire    [3:0]   i_ledlevel,
    input   wire    [1:0]   i_ledmode,
    input   wire    [1:0]   i_porta_status,
    input   wire    [1:0]   i_portb_status,
    input   wire    [1:0]   i_portc_status,
    input   wire    [1:0]   i_portd_status,
    input   wire    [11:0]  i_aio_dir,
    input   wire    [1:0]   i_harp_conf, // TODO
    input   wire    [15:0]  i_gpio_dir,  // TODO

    // Link power
    input   wire    [3:0]   i_link_pow,

    // HARP heartbeat
    input   wire            i_harp_hb,

    // Button press state
    input   wire    [5:0]   i_button,

    // Digital IO
    input   wire    [7:0]   i_din_state,
    input   wire    [7:0]   i_dout_state,

    // Neopixel control signal
    output  wire            o_neopix
);

//Timer for blinkenleds
parameter COUNTER_WIDTH = $clog2(CLK_RATE_HZ - 1);
reg [COUNTER_WIDTH - 1 : 0] counter = 'b0;
reg blink = 1'b1;

always @(posedge i_clk or posedge i_reset)
begin
    if (i_reset) begin
        counter <= 'b0;
        blink <= 1'b1;
    end else begin
        if (counter == CLK_RATE_HZ - 1) begin
            counter <= 'b0;
            blink <= ~blink;
        end else begin
            counter <= counter + 1'b1;
        end
    end
end

// Colors
reg [23:0] off,
           blue,
           orange,
           green,
           red,
           purple,
           brown ,
           pink ,
           white ,
           yellow,
           cyan;

// NB: This is hardcoded for the particular color set generated by colors.py
reg [23:0] colors [0:169];
reg [7:0] color_addr;
reg [3:0] color_idx, color_idx_last;
reg [23:0] color;

// Initialize RAM (produced by colors.py)
initial $readmemh("colors.mem", colors);
initial off = 0;

// RAM address
always @ (posedge i_clk) begin

    color_idx_last <= color_idx;

    if (i_reset) begin
        color_addr <= 0;
        color_idx <= 0;
    end else if (color_idx == 0) begin
        color_addr <= 153 + {4'b0000, i_ledlevel};
        color_idx <= 9;
    end else begin
        color_addr <= color_addr - 17;
        color_idx <= color_idx - 1;
    end
end

// RAM access
always @ (posedge i_clk) begin
    color <= colors[color_addr];
end

// Color update
always @ (posedge i_clk) begin
    case (color_idx_last)
        0: blue <= color;
        1: orange <= color;
        2: green <= color;
        3: red <= color;
        4: purple <= color;
        5: brown <= color;
        6: pink <= color;
        7: white <= color;
        8: yellow <= color;
        9: cyan <= color;
    endcase
end

// Neopixel color state
reg [23:0] rgb [0:40];

// LED on/off toggle 
reg dark = 1'b0;
reg [1:0] button0_history = 2'b00;

always @(posedge i_clk) begin

    button0_history <= {button0_history[0], i_button[0]};

    if (button0_history == 2'b01) begin
        dark <= dark + 1;
    end
end

// Port-specific running indicators
reg [3:0] port_running = 4'b0000;
reg [3:0] port_failed = 4'b0000;
reg last_acq_running = 1'b0;

always @(posedge i_clk) begin

    last_acq_running <= i_acq_running;

    // NB: Internal, port-specific running flag only changes on running start,
    // stop, or loss of lock or power
    if (!last_acq_running && i_acq_running) begin

        port_running <= {i_porta_status == 2'b11,
                         i_portb_status == 2'b11,
                         i_portc_status == 2'b11,
                         i_portd_status == 2'b11};
        port_failed <= 4'b0;

    end else if(!i_acq_running) begin

        port_running <= 4'b0;
        port_failed <= 4'b0;

    end else begin

        // Requires !i_acq_running to reset latch
        port_failed <= {port_failed[3] || (port_running[3] && i_porta_status != 2'b11),
                        port_failed[2] || (port_running[2] && i_portb_status != 2'b11),
                        port_failed[1] || (port_running[1] && i_portc_status != 2'b11),
                        port_failed[0] || (port_running[0] && i_portd_status != 2'b11)};
    end
end

wire leds_on = ~dark;

// LED color logic
always @(*) begin

    rgb[0] = leds_on ? yellow : off;

    rgb[1] = leds_on ?
            (i_acq_reset_done ?
            (i_acq_running ?
            (blink ?
            red : off) : red) : purple) : off;

    rgb[2] = (leds_on & i_button[5]) ? yellow : off;
    rgb[3] = (leds_on & i_button[4]) ? yellow : off;
    rgb[4] = (leds_on & i_button[3]) ? yellow : off;
    rgb[5] = (leds_on & i_button[2]) ? yellow : off;
    rgb[6] = (leds_on & i_button[1]) ? yellow : off;

    rgb[7] = (leds_on & i_harp_hb) ? red : off;
    rgb[8] = off; // TODO: "Host"

    rgb[9]  = (leds_on & i_dout_state[0]) ? blue : off;
    rgb[10] = (leds_on & i_dout_state[1]) ? blue : off;
    rgb[11] = (leds_on & i_dout_state[2]) ? blue : off;
    rgb[12] = (leds_on & i_dout_state[3]) ? blue : off;
    rgb[13] = (leds_on & i_dout_state[4]) ? blue : off;
    rgb[14] = (leds_on & i_dout_state[5]) ? blue : off;
    rgb[15] = (leds_on & i_dout_state[6]) ? blue : off;
    rgb[16] = (leds_on & i_dout_state[7]) ? blue : off;

    rgb[17] = (leds_on & i_din_state[7]) ? blue : off;
    rgb[18] = (leds_on & i_din_state[6]) ? blue : off;
    rgb[19] = (leds_on & i_din_state[5]) ? blue : off;
    rgb[20] = (leds_on & i_din_state[4]) ? blue : off;
    rgb[21] = (leds_on & i_din_state[3]) ? blue : off;
    rgb[22] = (leds_on & i_din_state[2]) ? blue : off;
    rgb[23] = (leds_on & i_din_state[1]) ? blue : off;
    rgb[24] = (leds_on & i_din_state[0]) ? blue : off;

    // NB: These if statements make heavy use of decending case priority
    // encoding

    // Port A (HS3 on the board)
    if (!leds_on || i_porta_status == 2'b00)            // Dark or power off
        rgb[25] = off;
    else if (port_failed[3])                            // Link issue in the middle of acquisition
        rgb[25] = orange;
    else if (port_running[3])                           // Acquisition running
        rgb[25] = blink ? red : off;
    else if (i_porta_status != 2'b01)                   // Locked
        rgb[25] = purple;
    else if (i_link_pow[3] && i_porta_status == 2'b01)  // Power on, waiting for lock
        rgb[25] = green;
    else
        rgb[25] = off;

    // Port B (HS2 on the board)
    if (!leds_on || i_portb_status == 2'b00)            // Dark or power off
        rgb[26] = off;
    else if (port_failed[2])                            // Link issue in the middle of acquisition
        rgb[26] = orange;
    else if (port_running[2])                           // Acquisition running
        rgb[26] = blink ? red : off;
    else if (i_portb_status != 2'b01)                   // Locked
        rgb[26] = purple;
    else if (i_link_pow[2] && i_portb_status == 2'b01)  // Power on, waiting for lock
        rgb[26] = green;
    else
        rgb[26] = off;

    // Port C (HS1 on the board)
    if (!leds_on || i_portc_status == 2'b00)            // Dark or power off
        rgb[27] = off;
    else if (port_failed[1])                            // Link issue in the middle of acquisition
        rgb[27] = orange;
    else if (port_running[1])                           // Acquisition running
        rgb[27] = blink ? red : off;
    else if (i_portc_status != 2'b01)                   // Locked
        rgb[27] = purple;
    else if (i_link_pow[1] && i_portc_status == 2'b01)  // Power on, waiting for lock
        rgb[27] = green;
    else
        rgb[27] = off;

    // Port D (HS0 on the board)
    if (!leds_on || i_portd_status == 2'b00)            // Dark or power off
        rgb[28] = off;
    else if (port_failed[0])                            // Link issue in the middle of acquisition
        rgb[28] = orange;
    else if (port_running[0])                           // Acquisition running
        rgb[28] = blink ? red : off;
    else if (i_portd_status != 2'b01)                   // Locked
        rgb[28] = purple;
    else if (i_link_pow[0] && i_portd_status == 2'b01)  // Power on, waiting for lock
        rgb[28] = green;
    else
        rgb[28] = off;

    // Analog IO. Input = green, output = red
    rgb[29] = leds_on ? (i_aio_dir[11] ? red : green) : off;
    rgb[30] = leds_on ? (i_aio_dir[10] ? red : green) : off;
    rgb[31] = leds_on ? (i_aio_dir[9]  ? red : green) : off;
    rgb[32] = leds_on ? (i_aio_dir[8]  ? red : green) : off;
    rgb[33] = leds_on ? (i_aio_dir[7]  ? red : green) : off;
    rgb[34] = leds_on ? (i_aio_dir[6]  ? red : green) : off;
    rgb[35] = leds_on ? (i_aio_dir[0]  ? red : green) : off;
    rgb[36] = leds_on ? (i_aio_dir[1]  ? red : green) : off;
    rgb[37] = leds_on ? (i_aio_dir[2]  ? red : green) : off;
    rgb[38] = leds_on ? (i_aio_dir[3]  ? red : green) : off;
    rgb[39] = leds_on ? (i_aio_dir[4]  ? red : green) : off;
    rgb[40] = leds_on ? (i_aio_dir[5]  ? red : green) : off;

end

// Currently addressed LED
wire [5:0] led_addr;

// Neopixel control
ws2811 # (
    .NUM_LEDS(41),
    .SYSTEM_CLOCK(CLK_RATE_HZ)
) neopix (
    .clk(i_clk),
    .reset(i_reset),
    .address(led_addr),
    .red_in(rgb[led_addr][23:16]),
    .green_in(rgb[led_addr][15:8]),
    .blue_in(rgb[led_addr][7:0]),
    .DO(o_neopix)
);

endmodule
